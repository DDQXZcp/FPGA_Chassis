//The following project is cotributed by Herman TANG
//No reproduction without permission.
module Top( 
	input ext_clk_50m,	//外部输入50MHz时钟信号
	input ext_rst_n,	//外部输入复位信号，低电平有效
////连接stm32
	input uart_rx,		// UART接收数据信号
	output uart_tx,		// UART发送数据信号			
//连接encoder
	input quadA,
	input quadB,
	output uart_clk,
	output quadA_test,
	output quadB_test,
	output uart_test,
	output total_pulse_test,
	output wire pwm0,pwm1,pwm2,pwm3
);

assign quadA_test = quadA;
assign quadB_test = quadB;	
//y_Global and X_Global are read directly from encoder, which is integer, one unit is related to physical configuration 
wire signed [31:0] y_Global,x_Global;

multiple_uart uart_controller (
    .clk(ext_clk_50m), 
    .rst_n(ext_rst_n), 
    .data1(x_Global[31:24]), //先用作测试
    .data2(x_Global[23:16]), 
    .data3(x_Global[15:8]), 
    .data4(x_Global[7:0]), 
    .uart_tx(uart_test), 
    .total_pulse_test(total_pulse_test)
    );
//return the 16bit encoder value						
quad Encoder_Y (
    .clk(ext_clk_50m), 
    .quadA(quadA), 
    .quadB(quadB), 
    .count(y_Global)
    );

quad Encoder_X (
    .clk(ext_clk_50m), 
    .quadA(quadA), 
    .quadB(quadB), 
    .count(x_Global)
    );

wire signed [31:0] current_x_speed;//current_Xspeed is derived from x_Global
wire signed [31:0] current_y_speed;//current_Xspeed is derived from y_Global
wire signed [31:0] current_angular_speed;//current_Xspeed is derived from y_Global
wire signed [31:0] target_x_speed;
wire signed [31:0] target_y_speed;
wire signed [31:0] target_angular_speed;
//need a speed calculation module

//The following setting is just for testing

assign target_x_speed = 32'd100000000;
assign target_y_speed = 32'd0;
assign target_angular_speed = 32'd0;//特殊说明：因为theta范围是0-65536

//need a module to generate target speed

wire [31:0] Kp,Ki,Kd;
assign Kp = 32'd4;//三位小数点
assign Ki = 32'd4;
assign Kd = 32'd4;
wire signed[39:0] x_speed, y_speed, angular_speed;// x_speed and y_speed is generated by PID controller

pid x_speed_pid (
    .clk(ext_clk_50m), 
    .nRst(ext_rst_n), 
    .target(target_x_speed), 
    .process(current_x_speed), 
    .Kp(Kp), 
    .Ki(Ki), 
    .Kd(Kd), 
    .drive(x_speed)
    );

pid y_speed_pid (
    .clk(ext_clk_50m), 
    .nRst(ext_rst_n), 
    .target(target_y_speed), 
    .process(current_y_speed), 
    .Kp(Kp), 
    .Ki(Ki), 
    .Kd(Kd), 
    .drive(y_speed)
    );

pid angular_speed_pid (
    .clk(ext_clk_50m), 
    .nRst(ext_rst_n), 
    .target(target_angular_speed), 
    .process(current_angular_speed), 
    .Kp(Kp), 
    .Ki(Ki), 
    .Kd(Kd), 
    .drive(angular_speed)
    );
	
//kinematic part

//theta preparation
wire [15:0] theta; //theta is unsigned, it can only range from 0-65536
theta_calculation theta_calculation (
    .clk(ext_clk_50m), 
    .rst_n(ext_rst_n), 
    .y_Global(y_Global), 
    .x_Global(x_Global), 
    .theta(theta)
    );
theta_calculation angular_speed_calculation (
    .clk(ext_clk_50m), 
    .rst_n(ext_rst_n), 
    .y_Global(current_x_speed), 
    .x_Global(current_x_speed), 
    .theta(current_angular_speed)
    );

// To test, if y_Global - x_Global is pi*L = 3.1415926*50 = 157, theta is 32768
wire signed[15:0] theta_sin,theta_cos;
wire signed[15:0] theta_sin_1,theta_cos_1;
wire signed[15:0] theta_sin_3,theta_cos_3;
wire signed[15:0] theta_sin_5,theta_cos_5;
wire signed[15:0] theta_sin_7,theta_cos_7;
//sin & cos value preparation
// -32767 represents -1.0 and +32767 represents +1.0.
//signed or unsigned for theta doesn't matter, the number is the same
//actually if no multiplication or division, no need to care the sign

//非常accurate, 使用isim进行仿真测试
icos theta_cos_converter1 (
    .x(theta), 
    .s(theta_cos)
    );
isin theta_sin_converter1 (
    .x(theta), 
    .s(theta_sin)
    );	
icos theta_cos_converter2 ( //pi = 32768, pi/4 = 8192
    .x(theta + 16'd8192), 
    .s(theta_cos_1)
    );
isin theta_sin_converter2 (
    .x(theta + 16'd8192), 
    .s(theta_sin_1)
    );	
icos theta_cos_converter3 ( //pi = 32768, pi*3/4 = 24576
    .x(theta + 16'd24576), 
    .s(theta_cos_3)
    );
isin theta_sin_converter3 (
    .x(theta + 16'd24576), 
    .s(theta_sin_3)
    );	
icos theta_cos_converter4 ( //pi = 32768, pi*3/4 = 24576
    .x(theta - 16'd24576), 
    .s(theta_cos_5)
    );
isin theta_sin_converter4 (
    .x(theta - 16'd24576), 
    .s(theta_sin_5)
    );	
icos theta_cos_converter5 ( //pi = 32768, pi*3/4 = 24576
    .x(theta - 16'd8192), 
    .s(theta_cos_7)
    );
isin theta_sin_converter5 (
    .x(theta - 16'd8192), 
    .s(theta_sin_7)
    );	

//kinematic calculation
//To convert the desired global speed to the speed of each motor
// pi = 65536/2 = 32768,theta is 16bit
/*  The C program
	Rspeed[0] = Gvx * (-1) * sin(theta + pi / 4) + Gvy * cos(theta + pi / 4) + r * theta;
    Rspeed[1] = Gvx * (-1) * sin(theta + 3 * pi / 4) + Gvy * cos(theta + 3 * pi / 4) + r * theta;
    Rspeed[2] = Gvx * (-1) * sin(theta + 5 * pi / 4) + Gvy * cos(theta + 5 * pi / 4) + r * theta;
    Rspeed[3] = Gvx * (-1) * sin(theta + 7 * pi / 4) + Gvy * cos(theta + 7 * pi / 4) + r * theta;
*/
wire signed[55:0] MotorSpeed0,MotorSpeed1,MotorSpeed2,MotorSpeed3;
// Take care the range theta_cos_x and theta_sin_x range from -32767 ~ 32767
//The result is scaled to 2^15 2^16?
parameter L = 50;// This L is the distance from motor to the center of chassis
//MotorSpeed -32767~32767 is multiplied by a scale of -32767~32767, become a 32-bit data
//y_speed 40 bit, theta_cos 16 bit
assign	MotorSpeed0 = y_speed * theta_cos_1 - x_speed * theta_sin_1 + L * angular_speed; 
assign	MotorSpeed1 = y_speed * theta_cos_3 - x_speed * theta_sin_3 + L * angular_speed;
assign	MotorSpeed2 = y_speed * theta_cos_5 - x_speed * theta_sin_5 + L * angular_speed; 
assign	MotorSpeed3 = y_speed * theta_cos_7 - x_speed * theta_sin_7 + L * angular_speed; 

// DC motor pwm control, 16 bit resolution
//need to convert the signed to unsigned
//Check the signed bit, if signed, do 2's complement and control the H bridge
wire Hbridge1,Hbridge2;
wire Hbridge3,Hbridge4;
wire Hbridge5,Hbridge6;
wire Hbridge7,Hbridge8;
pwmmodule motor_pwm_output0 (
    .data(MotorSpeed0[55:16]),//automatically divided by 2^16
    .reset(ext_rst_n), 
    .clk(ext_clk_50m), 
    .pwm(pwm0), 
    .Hbridge1(Hbridge1), 
    .Hbridge2(Hbridge2)
    );
pwmmodule motor_pwm_output1 (
    .data(MotorSpeed1[55:16]),//automatically divided by 2^16
    .reset(ext_rst_n), 
    .clk(ext_clk_50m), 
    .pwm(pwm1), 
    .Hbridge1(Hbridge3), 
    .Hbridge2(Hbridge4)
    );
pwmmodule motor_pwm_output2 (
    .data(MotorSpeed2[55:16]),//automatically divided by 2^16
    .reset(ext_rst_n), 
    .clk(ext_clk_50m), 
    .pwm(pwm2), 
    .Hbridge1(Hbridge5), 
    .Hbridge2(Hbridge6)
    );
pwmmodule motor_pwm_output3 (
    .data(MotorSpeed3[55:16]),//automatically divided by 2^16
    .reset(ext_rst_n), 
    .clk(ext_clk_50m), 
    .pwm(pwm3), 
    .Hbridge1(Hbridge7), 
    .Hbridge2(Hbridge8)
    );


endmodule